module MemInstrucoes ( adress , Instrucao , clock, clockAUTO ) ;

 input [9:0] adress ;
 input clockAUTO;
 input clock ;
 output [31:0] Instrucao ;
 reg [31:0] mem [255:0];
 integer flag = 0;
 
 reg[31:0] x;

 always @ ( negedge clock )
 begin
 if ( flag == 0)
 begin
 // PAR OU IMPAR
 /*
 mem[0] =  32'b01101100000000000000000000000000;  //nop
 mem[1] =  32'b01011100001000000000000000000000;  //in
 mem[2] =  32'b01000000000000100000000000000010; // r[2] = 2;
 mem[3] =  32'b01100100010000100000000000000101; // r[2] = r[2] << 5;
 mem[4] =  32'b01101000010000100000000000000101; // r[2] = r[2] >> 5;
 mem[5] =  32'b00010000001000100001100000000000; // r[3] = r[1] % r[2];
 mem[6] =  32'b00011100011000000000000000001010; // bgt r[3] > r[0], PC=10
 mem[10] =  32'b00100000000000110000000000001100; // blt r[0] > r[3], PC=12
 mem[12] =  32'b00101100011000000000000000001110; // bgtz r[3] > 0, PC=14
 mem[14] =  32'b01100000011000000000000000000000;  //out
 mem[15] =  32'b01110000000000000000000000000000;  //halt
 */
 
 //TESTE XOR
 /*
 mem[0] =  32'b01101100000000000000000000000000;  //nop
 mem[1] =  32'b01011100000000000000000000000000;  //in
 mem[2] =  32'b01001100001000100000000000000100; // slti r[2], r[1] < 4
 mem[3] =  32'b00010100000000100000000000000101; // beq r[2] == r[0], PC=5
 mem[4] =  32'b01011000001000010000100000000000; //r1 = r1 xor r1
 mem[5] =  32'b01100000001000000000000000000000;  //out
 mem[6] =  32'b01110000000000000000000000000000;  //halt
 */

 
 //FIBONACCI 1
 /*
 mem[0] =  32'b01101100000000000000000000000000;  //nop
 mem[1] =  32'b01011100000000000000000000000000;  //in
 mem[2] =  32'b00001100001000100000000000000001;  //r[2]=r[1]-1
 mem[3] =  32'b01000000000001010000000000000001; // r[5] = 1;
 mem[5] =  32'b01000000000000110000000000000000; // r[3] = 0;
 mem[6] =  32'b010000/00000/00100/0000000000000001; // r[4] = 1;
 mem[7] =  32'b01001000000000100101000000000000; // slt r[10], r[0], r[2]
 mem[8] =  32'b00010100000010100000000000010001; // beq r[10] == r[0], PC=17
 mem[9] =  32'b00011000000010100000000000001010; // bne r[10] != r[0], PC=10
 mem[10] = 32'b00000000011001000010100000000000; //r5 = r3 + r4
 mem[11] = 32'b01010100101000000010100000000000; //r5 = r5 ou r0
 mem[12] = 32'b00000000100000000001100000000000; //r3 = r4
 mem[13] = 32'b00000000101000000010000000000000; //r4 = r5
 mem[14] = 32'b00001100010000100000000000000001;  //r[2]=r[2]-1
 mem[15] = 32'b00110100000000000000000000000111;  //pc=7
 mem[16] = 32'b01010000101000000010100000000000; //r5 = r5 and r0
 mem[17] = 32'b01100000101000000000000000000000;  //out
 mem[18] = 32'b01110000000000000000000000000000;  //halt 
 */
 
 
 
 //FATORIAL
 /*
 mem[0] =  32'b01101100000000000000000000000000;  //nop
 mem[1] =  32'b010111_00001_000000000000000000000;  //in
 mem[2] =  32'b00001100001000100000000000000001;  //r[2]=r[1]-1
 mem[3] =  32'b01001000000000100101000000000000; // slt r[10], r[0], r[2]
 mem[4] =  32'b00010100000010100000000000001000; // beq r[10] == r[0], PC=8
 mem[5] =  32'b00110000001000100000100000000000;  //r[1] = r[1]*r[2]
 mem[6] =  32'b00001100010000100000000000000001;  //r[2]=r[2]-1
 mem[7] =  32'b00110100000000000000000000000011;  //pc=3
 mem[8] =  32'b01100000001000000000000000000010;  //out
 mem[9] =  32'b01110000000000000000000000000000;  //halt
 */
 
	//SELECTION
	/*
	mem[0]	=	32'b010000_00000_11011_0000000000000000;
	mem[1]	=	32'b010000_00000_11100_0000000000101000;
	mem[2]	=	32'b010000_00000_11101_0000000000110010;
	mem[3]	=	32'b001101_00000000000000000001111101;
	mem[4]	=	32'b010001_11011_10001_0000000000000000;
	mem[5]	=	32'b010001_11011_10010_0000000000000001;
	mem[6]	=	32'b010001_11011_10011_0000000000000010;
	mem[7]	=	32'b001111_11011_00001_0000000000000101;
	mem[8]	=	32'b001111_11011_00010_0000000000000001;
	mem[9]	=	32'b011101_00010_00001_0000000000000000;
	mem[10]	=	32'b010001_11011_00001_0000000000000101;
	mem[11]	=	32'b001111_11011_00011_0000000000000100;
	mem[12]	=	32'b001111_11011_00101_0000000000000001;
	mem[13]	=	32'b001111_11011_00100_0000000000000000;
	mem[14]	=	32'b000000_00101_00100_00101_00000000000;
	mem[15]	=	32'b001111_00101_00100_0000000000000000;
	mem[16]	=	32'b011101_00100_00011_0000000000000000;
	mem[17]	=	32'b010001_11011_00011_0000000000000100;
	mem[18]	=	32'b001111_11011_00110_0000000000000011;
	mem[19]	=	32'b001111_11011_00111_0000000000000001;
	mem[20]	=	32'b010000_00000_01000_0000000000000001;
	mem[21]	=	32'b000000_00111_01000_01001_00000000000;
	mem[22]	=	32'b011101_01001_00110_0000000000000000;
	mem[23]	=	32'b010001_11011_00110_0000000000000011;
	mem[24]	=	32'b001111_11011_01010_0000000000000011;
	mem[25]	=	32'b001111_11011_01011_0000000000000010;
	mem[26]	=	32'b010010_01010_01011_01100_00000000000;
	mem[27]	=	32'b000101_01100_00000_0000000000110110;
	mem[28]	=	32'b001111_11011_01110_0000000000000011;
	mem[29]	=	32'b001111_11011_01101_0000000000000000;
	mem[30]	=	32'b000000_01110_01101_01110_00000000000;
	mem[31]	=	32'b001111_01110_01101_0000000000000000;
	mem[32]	=	32'b001111_11011_01111_0000000000000100;
	mem[33]	=	32'b010010_01101_01111_10000_00000000000;
	mem[34]	=	32'b000101_10000_00000_0000000000101111;
	mem[35]	=	32'b001111_11011_00001_0000000000000100;
	mem[36]	=	32'b001111_11011_00011_0000000000000011;
	mem[37]	=	32'b001111_11011_00010_0000000000000000;
	mem[38]	=	32'b000000_00011_00010_00011_00000000000;
	mem[39]	=	32'b001111_00011_00010_0000000000000000;
	mem[40]	=	32'b011101_00010_00001_0000000000000000;
	mem[41]	=	32'b010001_11011_00001_0000000000000100;
	mem[42]	=	32'b001111_11011_00100_0000000000000101;
	mem[43]	=	32'b001111_11011_00101_0000000000000011;
	mem[44]	=	32'b011101_00101_00100_0000000000000000;
	mem[45]	=	32'b010001_11011_00100_0000000000000101;
	mem[46]	=	32'b001101_00000000000000000000101111;
	mem[47]	=	32'b001111_11011_00110_0000000000000011;
	mem[48]	=	32'b001111_11011_00111_0000000000000011;
	mem[49]	=	32'b010000_00000_01000_0000000000000001;
	mem[50]	=	32'b000000_00111_01000_01001_00000000000;
	mem[51]	=	32'b011101_01001_00110_0000000000000000;
	mem[52]	=	32'b010001_11011_00110_0000000000000011;
	mem[53]	=	32'b001101_00000000000000000000011000;
	mem[54]	=	32'b001111_11011_01010_0000000000000101;
	mem[55]	=	32'b011101_01010_11110_0000000000000000;
	mem[56]	=	32'b000001_11101_11101_1111111111111111;
	mem[57]	=	32'b001111_11101_11111_0000000000000000;
	mem[58]	=	32'b001110_11111_00000_0000000000000000;
	mem[59]	=	32'b000001_11101_11101_1111111111111111;
	mem[60]	=	32'b001111_11101_11111_0000000000000000;
	mem[61]	=	32'b001110_11111_00000_0000000000000000;
	mem[62]	=	32'b010001_11011_10001_0000000000000000;
	mem[63]	=	32'b010001_11011_10010_0000000000000001;
	mem[64]	=	32'b010001_11011_10011_0000000000000010;
	mem[65]	=	32'b001111_11011_01011_0000000000000011;
	mem[66]	=	32'b001111_11011_01100_0000000000000001;
	mem[67]	=	32'b011101_01100_01011_0000000000000000;
	mem[68]	=	32'b010001_11011_01011_0000000000000011;
	mem[69]	=	32'b001111_11011_01101_0000000000000011;
	mem[70]	=	32'b001111_11011_01110_0000000000000010;
	mem[71]	=	32'b010000_00000_01111_0000000000000001;
	mem[72]	=	32'b000010_01110_01111_10000_00000000000;
	mem[73]	=	32'b010010_01101_10000_00001_00000000000;
	mem[74]	=	32'b000101_00001_00000_0000000001111010;
	mem[75]	=	32'b001111_11011_00010_0000000000000100;
	mem[76]	=	32'b001111_11011_00011_0000000000000000;
	mem[77]	=	32'b011101_00011_10001_0000000000000000;
	mem[78]	=	32'b001111_11011_00100_0000000000000011;
	mem[79]	=	32'b011101_00100_10010_0000000000000000;
	mem[80]	=	32'b001111_11011_00101_0000000000000010;
	mem[81]	=	32'b011101_00101_10011_0000000000000000;
	mem[82]	=	32'b000001_11011_11011_0000000000000110;
	mem[83]	=	32'b010000_00000_11111_0000000001010111;
	mem[84]	=	32'b010001_11101_11111_0000000000000000;
	mem[85]	=	32'b000001_11101_11101_0000000000000001;
	mem[86]	=	32'b001101_00000000000000000000000100;
	mem[87]	=	32'b011101_11110_00110_0000000000000000;
	mem[88]	=	32'b000001_11011_11011_1111111111111010;
	mem[89]	=	32'b011101_00110_00010_0000000000000000;
	mem[90]	=	32'b010001_11011_00010_0000000000000100;
	mem[91]	=	32'b001111_11011_00111_0000000000000101;
	mem[92]	=	32'b001111_11011_01001_0000000000000100;
	mem[93]	=	32'b001111_11011_01000_0000000000000000;
	mem[94]	=	32'b000000_01001_01000_01001_00000000000;
	mem[95]	=	32'b001111_01001_01000_0000000000000000;
	mem[96]	=	32'b011101_01000_00111_0000000000000000;
	mem[97]	=	32'b010001_11011_00111_0000000000000101;
	mem[98]	=	32'b001111_11011_01011_0000000000000100;
	mem[99]	=	32'b001111_11011_01010_0000000000000000;
	mem[100]	=	32'b000000_01011_01010_01011_00000000000;
	mem[101]	=	32'b001111_01011_01010_0000000000000000;
	mem[102]	=	32'b001111_11011_01101_0000000000000011;
	mem[103]	=	32'b001111_11011_01100_0000000000000000;
	mem[104]	=	32'b000000_01101_01100_01101_00000000000;
	mem[105]	=	32'b001111_01101_01100_0000000000000000;
	mem[106]	=	32'b011101_01100_01010_0000000000000000;
	mem[107]	=	32'b010001_01011_01010_0000000000000000;
	mem[108]	=	32'b001111_11011_01111_0000000000000011;
	mem[109]	=	32'b001111_11011_01110_0000000000000000;
	mem[110]	=	32'b000000_01111_01110_01111_00000000000;
	mem[111]	=	32'b001111_01111_01110_0000000000000000;
	mem[112]	=	32'b001111_11011_10000_0000000000000101;
	mem[113]	=	32'b011101_10000_01110_0000000000000000;
	mem[114]	=	32'b010001_01111_01110_0000000000000000;
	mem[115]	=	32'b001111_11011_00001_0000000000000011;
	mem[116]	=	32'b001111_11011_00010_0000000000000011;
	mem[117]	=	32'b010000_00000_00011_0000000000000001;
	mem[118]	=	32'b000000_00010_00011_00100_00000000000;
	mem[119]	=	32'b011101_00100_00001_0000000000000000;
	mem[120]	=	32'b010001_11011_00001_0000000000000011;
	mem[121]	=	32'b001101_00000000000000000001000101;
	mem[122]	=	32'b000001_11101_11101_1111111111111111;
	mem[123]	=	32'b001111_11101_11111_0000000000000000;
	mem[124]	=	32'b001110_11111_00000_0000000000000000;
	mem[125]	=	32'b001111_11011_00101_0000000000000000;
	mem[126]	=	32'b010000_00000_00110_0000000000000000;
	mem[127]	=	32'b011101_00110_00101_0000000000000000;
	mem[128]	=	32'b010001_11011_00101_0000000000000000;
	mem[129]	=	32'b001111_11011_00111_0000000000000000;
	mem[130]	=	32'b010000_00000_01000_0000000000000011;
	mem[131]	=	32'b010010_00111_01000_01001_00000000000;
	mem[132]	=	32'b000101_01001_00000_0000000010010010;
	mem[133]	=	32'b001111_11011_01011_0000000000000000;
	mem[134]	=	32'b000000_01011_11100_01011_00000000000;
	mem[135]	=	32'b001111_01011_01010_0000000000000000;
	mem[136]	=	32'b010111_01100_00000_0000000000000000;
	mem[137]	=	32'b011101_01100_01010_0000000000000000;
	mem[138]	=	32'b010001_01011_01010_0000000000000000;
	mem[139]	=	32'b001111_11011_01101_0000000000000000;
	mem[140]	=	32'b001111_11011_01110_0000000000000000;
	mem[141]	=	32'b010000_00000_01111_0000000000000001;
	mem[142]	=	32'b000000_01110_01111_10000_00000000000;
	mem[143]	=	32'b011101_10000_01101_0000000000000000;
	mem[144]	=	32'b010001_11011_01101_0000000000000000;
	mem[145]	=	32'b001101_00000000000000000010000001;
	mem[146]	=	32'b000001_11100_00001_0000000000000000;
	mem[147]	=	32'b011101_00001_10001_0000000000000000;
	mem[148]	=	32'b010000_00000_00010_0000000000000000;
	mem[149]	=	32'b011101_00010_10010_0000000000000000;
	mem[150]	=	32'b010000_00000_00011_0000000000000011;
	mem[151]	=	32'b011101_00011_10011_0000000000000000;
	mem[152]	=	32'b000001_11011_11011_0000000000000001;
	mem[153]	=	32'b010000_00000_11111_0000000010011101;
	mem[154]	=	32'b010001_11101_11111_0000000000000000;
	mem[155]	=	32'b000001_11101_11101_0000000000000001;
	mem[156]	=	32'b001101_00000000000000000000111110;
	mem[157]	=	32'b011101_11110_00100_0000000000000000;
	mem[158]	=	32'b000001_11011_11011_1111111111111111;
	mem[159]	=	32'b001111_11011_00101_0000000000000000;
	mem[160]	=	32'b010000_00000_00110_0000000000000000;
	mem[161]	=	32'b011101_00110_00101_0000000000000000;
	mem[162]	=	32'b010001_11011_00101_0000000000000000;
	mem[163]	=	32'b001111_11011_00111_0000000000000000;
	mem[164]	=	32'b010000_00000_01000_0000000000000011;
	mem[165]	=	32'b010010_00111_01000_01001_00000000000;
	mem[166]	=	32'b000101_01001_00000_0000000010110101;
	mem[167]	=	32'b001111_11011_01011_0000000000000000;
	mem[168]	=	32'b000000_01011_11100_01011_00000000000;
	mem[169]	=	32'b001111_01011_01010_0000000000000000;
	mem[170]	=	32'b011101_01010_10001_0000000000000000;
	mem[171]	=	32'b011101_10001_01100_0000000000000000;
	mem[172]	=	32'b011000_01100_00000_0000000000000000;
	mem[173]	=	32'b011011_00000000000000000000000000;
	mem[174]	=	32'b001111_11011_01101_0000000000000000;
	mem[175]	=	32'b001111_11011_01110_0000000000000000;
	mem[176]	=	32'b010000_00000_01111_0000000000000001;
	mem[177]	=	32'b000000_01110_01111_10000_00000000000;
	mem[178]	=	32'b011101_10000_01101_0000000000000000;
	mem[179]	=	32'b010001_11011_01101_0000000000000000;
	mem[180]	=	32'b001101_00000000000000000010100011;
	mem[181]	=	32'b001101_00000000000000000010110110;
	mem[182]	=	32'b011100_00000000000000000000000000;
	*/
	
	//GCD
	
	mem[0]	=	32'b010000_00000_11011_0000000000000000;
	mem[1]	=	32'b010000_00000_11100_0000000000101000;
	mem[2]	=	32'b010000_00000_11101_0000000000110010;
	mem[3]	=	32'b001101_00000000000000000000101011;
	mem[4]	=	32'b010001_11011_10001_0000000000000000;
	mem[5]	=	32'b010001_11011_10010_0000000000000001;
	mem[6]	=	32'b001111_11011_00001_0000000000000001;
	mem[7]	=	32'b010000_00000_00010_0000000000000000;
	mem[8]	=	32'b100000_00001_00010_00011_00000000000;
	mem[9]	=	32'b011111_00001_00010_00100_00000000000;
	mem[10]	=	32'b010100_00011_00100_00101_00000000000;
	mem[11]	=	32'b000101_00101_00000_0000000000010010;
	mem[12]	=	32'b001111_11011_00110_0000000000000000;
	mem[13]	=	32'b011101_00110_11110_0000000000000000;
	mem[14]	=	32'b000001_11101_11101_1111111111111111;
	mem[15]	=	32'b001111_11101_11111_0000000000000000;
	mem[16]	=	32'b001110_11111_00000_0000000000000000;
	mem[17]	=	32'b001101_00000000000000000000101000;
	mem[18]	=	32'b001111_11011_00111_0000000000000001;
	mem[19]	=	32'b011101_00111_10001_0000000000000000;
	mem[20]	=	32'b001111_11011_01000_0000000000000000;
	mem[21]	=	32'b001111_11011_01001_0000000000000000;
	mem[22]	=	32'b001111_11011_01010_0000000000000001;
	mem[23]	=	32'b100001_01001_01010_01011_00000000000;
	mem[24]	=	32'b001111_11011_01100_0000000000000001;
	mem[25]	=	32'b001100_01011_01100_01101_00000000000;
	mem[26]	=	32'b000010_01000_01101_01110_00000000000;
	mem[27]	=	32'b011101_01110_10010_0000000000000000;
	mem[28]	=	32'b000001_11011_11011_0000000000000010;
	mem[29]	=	32'b010000_00000_11111_0000000000100001;
	mem[30]	=	32'b010001_11101_11111_0000000000000000;
	mem[31]	=	32'b000001_11101_11101_0000000000000001;
	mem[32]	=	32'b001101_00000000000000000000000100;
	mem[33]	=	32'b011101_11110_01111_0000000000000000;
	mem[34]	=	32'b000001_11011_11011_1111111111111110;
	mem[35]	=	32'b011101_01111_11110_0000000000000000;
	mem[36]	=	32'b000001_11101_11101_1111111111111111;
	mem[37]	=	32'b001111_11101_11111_0000000000000000;
	mem[38]	=	32'b001110_11111_00000_0000000000000000;
	mem[39]	=	32'b001101_00000000000000000000101000;
	mem[40]	=	32'b000001_11101_11101_1111111111111111;
	mem[41]	=	32'b001111_11101_11111_0000000000000000;
	mem[42]	=	32'b001110_11111_00000_0000000000000000;
	mem[43]	=	32'b001111_11011_10000_0000000000000000;
	mem[44]	=	32'b010111_00001_00000_0000000000000000;
	mem[45]	=	32'b011101_00001_10000_0000000000000000;
	mem[46]	=	32'b010001_11011_10000_0000000000000000;
	mem[47]	=	32'b001111_11011_00010_0000000000000001;
	mem[48]	=	32'b010111_00011_00000_0000000000000000;
	mem[49]	=	32'b011101_00011_00010_0000000000000000;
	mem[50]	=	32'b010001_11011_00010_0000000000000001;
	mem[51]	=	32'b001111_11011_00100_0000000000000000;
	mem[52]	=	32'b011101_00100_10001_0000000000000000;
	mem[53]	=	32'b001111_11011_00101_0000000000000001;
	mem[54]	=	32'b011101_00101_10010_0000000000000000;
	mem[55]	=	32'b000001_11011_11011_0000000000000010;
	mem[56]	=	32'b010000_00000_11111_0000000000111100;
	mem[57]	=	32'b010001_11101_11111_0000000000000000;
	mem[58]	=	32'b000001_11101_11101_0000000000000001;
	mem[59]	=	32'b001101_00000000000000000000000100;
	mem[60]	=	32'b011101_11110_00110_0000000000000000;
	mem[61]	=	32'b000001_11011_11011_1111111111111110;
	mem[62]	=	32'b011101_00110_10001_0000000000000000;
	mem[63]	=	32'b011101_10001_00111_0000000000000000;
	mem[64]	=	32'b011000_00111_00000_0000000000000000;
	mem[65]	=	32'b011011_00000000000000000000000000;
	mem[66]	=	32'b001101_00000000000000000001000011;
	mem[67]	=	32'b011100_00000000000000000000000000;
	




	
 //FIBONACCI 2
 /*
 mem[0] =  32'b01101100000000000000000000000000;  //nop
 mem[1] =  32'b01011100001000000000000000000000;  //in
 mem[2] =  32'b00001100001000100000000000000001;  //r[2]=r[1]-1
 mem[3] =  32'b01000000000001100000000000001001; // r[6] = 9;
 mem[4] =  32'b01000000000010110000000000000001; // r[11] = 1;
 mem[5] =  32'b01000000000001010000000000000001; // r[5] = 1;
 mem[6] =  32'b01000000000000110000000000000000; // r[3] = 0;
 mem[7] =  32'b01000100000001010000000000000001; // m[1] = r[5]
 mem[8] =  32'b00111100000001000000000000000001; // r[4] = m[1];
 mem[9] =  32'b01001000000000100101000000000000; // slt r[10], r[0], r[2]
 mem[10] = 32'b00100100000010100000000000010001; // beqz r[10] == 0, PC=17
 mem[11] = 32'b00101000000010100000000000001100; // bnez r[10] != 0, PC=12
 mem[12] = 32'b00000000011001000010100000000000; //r5 = r3 + r4
 mem[13] = 32'b00000000100000000001100000000000; //r3 = r4
 mem[14] = 32'b00000000101000000010000000000000; //r4 = r5
 mem[15] = 32'b00001000010010110001000000000000;  //r[2]=r[2]-r[11]
 mem[16] = 32'b00111000110000000000000000000000;  //pc=r[6]
 mem[17] = 32'b01100000101000000000000000000010;  //out
 mem[18] =  32'b01110000000000000000000000000000;  //halt 
 
 */
 

 
 

 
flag <= 1;
 end
 end
 
 always @ ( negedge clockAUTO )
 begin
 x <= mem [ adress ];
 end
 
 assign Instrucao = x;
 endmodule
