module display_verilog(entrada, clock_atual, saida1,saida2,saida3,saida4,saida_clock1,saida_clock2,traco);

	input [31:0] entrada;
	input [9:0] clock_atual;
	output reg[6:0]saida1;
	output reg[6:0]saida2;
	output reg[6:0]saida3;
	output reg[6:0]saida4;
	output reg[6:0]saida_clock1;
	output reg[6:0]saida_clock2;
	output reg[1:0]traco;
	reg [31:0] d1;
	reg [31:0] d2;
	reg [31:0] d3;
	reg [31:0] d4;
	reg [31:0] c1;
	reg [31:0] c2;
	
	always@(*)
	
		begin	
		
		traco = 2'b00;
		
			if(entrada < 10)
				begin
			
				saida2 = 7'b0000001;
				saida3 = 7'b0000001;
				saida4 = 7'b0000001;
				
				case (entrada)
				
					32'b00000000000000000000000000000000: saida1 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida1 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida1 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida1 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida1 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida1 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida1 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida1 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida1 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida1 = 7'b0000100;
				
				endcase	
				end
			
			
			else if((entrada>=10) && (entrada<100)) 
				
				begin
			
				d1 = entrada % 10;
				d2 = entrada / 10;
				saida3 = 7'b0000001;
				saida4 = 7'b0000001;
				
				case (d1)
				
					32'b00000000000000000000000000000000: saida1 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida1 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida1 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida1 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida1 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida1 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida1 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida1 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida1 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida1 = 7'b0000100;
				
			
			endcase
			
			case (d2)
				
					32'b00000000000000000000000000000000: saida2 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida2 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida2 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida2 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida2 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida2 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida2 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida2 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida2 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida2 = 7'b0000100;
				
				endcase
			end
			
			else if((entrada>=100) && (entrada<1000))
			
				begin
			
				d1 = entrada % 100;
				d1 = d1 % 10;
				d2 = entrada / 10;
				d2 = d2 % 10;
				d3 = entrada / 100;
				saida4 = 7'b0000001;
				
				case (d1)
				
					32'b00000000000000000000000000000000: saida1 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida1 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida1 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida1 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida1 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida1 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida1 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida1 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida1 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida1 = 7'b0000100;
				
			
			endcase
			
			case (d2)
				
					32'b00000000000000000000000000000000: saida2 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida2 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida2 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida2 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida2 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida2 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida2 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida2 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida2 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida2 = 7'b0000100;
				
				endcase
				
			case (d3)
				
					32'b00000000000000000000000000000000: saida3 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida3 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida3 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida3 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida3 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida3 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida3 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida3 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida3 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida3 = 7'b0000100;
				
				endcase
			end
	
		else if(entrada>=1000)
			
				begin
			
				d1 = entrada % 10;
				d2 = entrada / 10;
				d2 = d2 % 10;
				d3 = entrada / 100;
				d3 = d3 % 10;
				d4 = entrada / 1000;
				
				case (d1)
				
					32'b00000000000000000000000000000000: saida1 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida1 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida1 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida1 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida1 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida1 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida1 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida1 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida1 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida1 = 7'b0000100;
				
			
			endcase
			
			case (d2)
				
					32'b00000000000000000000000000000000: saida2 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida2 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida2 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida2 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida2 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida2 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida2 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida2 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida2 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida2 = 7'b0000100;
				
				endcase
				
			case (d3)
				
					32'b00000000000000000000000000000000: saida3 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida3 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida3 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida3 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida3 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida3 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida3 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida3 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida3 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida3 = 7'b0000100;
				
				endcase
				
			case (d4)
				
					32'b00000000000000000000000000000000: saida4 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida4 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida4 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida4 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida4 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida4 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida4 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida4 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida4 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida4 = 7'b0000100;
				
				endcase
			end
			
		end
	
	
	
	
	always@(clock_atual)
			
			begin
			
			if(clock_atual<10)
			
			begin
			
			saida_clock2 = 7'b0000001;
			
			case (clock_atual)
				
					32'b00000000000000000000000000000000: saida_clock1 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida_clock1 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida_clock1 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida_clock1 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida_clock1 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida_clock1 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida_clock1 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida_clock1 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida_clock1 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida_clock1 = 7'b0000100;
				
				endcase
			end
			
			else if(clock_atual>=10)
			
			begin
			
			c1 = clock_atual % 10;
			c2 = clock_atual/10;
			
			case (c1)
				
					32'b00000000000000000000000000000000: saida_clock1 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida_clock1 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida_clock1 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida_clock1 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida_clock1 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida_clock1 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida_clock1 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida_clock1 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida_clock1 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida_clock1 = 7'b0000100;
				
				endcase
				
			case (c2)
				
					32'b00000000000000000000000000000000: saida_clock2 = 7'b0000001; 
					32'b00000000000000000000000000000001: saida_clock2 = 7'b1001111; 
					32'b00000000000000000000000000000010: saida_clock2 = 7'b0010010; 
					32'b00000000000000000000000000000011: saida_clock2 = 7'b0000110; 
					32'b00000000000000000000000000000100: saida_clock2 = 7'b1001100; 
					32'b00000000000000000000000000000101: saida_clock2 = 7'b0100100; 
					32'b00000000000000000000000000000110: saida_clock2 = 7'b0100000; 
					32'b00000000000000000000000000000111: saida_clock2 = 7'b0001111; 
					32'b00000000000000000000000000001000: saida_clock2 = 7'b0000000; 
					32'b00000000000000000000000000001001: saida_clock2 = 7'b0000100;
				
				endcase
			end
		end
	

	endmodule

