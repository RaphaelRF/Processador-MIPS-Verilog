module Input (data,in, clock,saida);

input [3:0] data;
input clock, in;
output reg [31:0] saida;

always @ ( posedge clock )
begin
if(in)

case(data)

4'b0000: saida = 32'b00000000000000000000000000000000;
4'b0001: saida = 32'b00000000000000000000000000000001;
4'b0010: saida = 32'b00000000000000000000000000000010;
4'b0011: saida = 32'b00000000000000000000000000000011;
4'b0100: saida = 32'b00000000000000000000000000000100;
4'b0101: saida = 32'b00000000000000000000000000000101;
4'b0110: saida = 32'b00000000000000000000000000000110;
4'b0111: saida = 32'b00000000000000000000000000000111;
4'b1000: saida = 32'b00000000000000000000000000001000;
4'b1001: saida = 32'b00000000000000000000000000001001;
4'b1010: saida = 32'b00000000000000000000000000001010;
4'b1011: saida = 32'b00000000000000000000000000001011;
4'b1100: saida = 32'b00000000000000000000000000001100;
4'b1101: saida = 32'b00000000000000000000000000001101;
4'b1110: saida = 32'b00000000000000000000000000001110;
4'b1111: saida = 32'b00000000000000000000000000001111;
//3'b111: saida = 32'b00000000000000000000000000000000;
default saida = 32'b00000000000000000000000000000000;
endcase
end

endmodule
